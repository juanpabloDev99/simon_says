library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity buttonsInterface_tb is
end buttonsInterface_tb;

architecture Behavioral of buttonsInterface_tb is

begin

end Behavioral;
